// Description: Common RISC-V definitions

package riscv;

    localparam VLEN = 32; //virtual address length
    localparam PLEN = 34; //physical address length

endpackage
